////////////////////////////////////////////////////////////////////////////////
// Adder
////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps 

module Adder(
    input [3:0] a,b,
    output [3:0] c
);

    assign c = a+b;
    
endmodule
