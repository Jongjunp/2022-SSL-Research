`timescale 1ns / 1ps 

module tester #(
    parameter A = 8,
    parameter B = 8,
    parameter ADDER_0 = A + 1
)
(
    input wire                  ;
    input 
);

    initial
    begin



    end
    